`timescale 1 ns / 1ps

module InstrMem (
    input [31:0] cur_pc,
    output reg [31:0] instruction
);

    reg [7:0] rom[311:0];
    integer i;

// initialization
    initial begin
        for(i=0;i<511;i=i+1)begin
            rom[i] = 8'b0000_0000;
        end
        {rom[3],rom[2],rom[1],rom[0]} = 32'b00011001001100000000001010010011;
        {rom[7],rom[6],rom[5],rom[4]} = 32'b00000000000000000000000000010011;
        {rom[11],rom[10],rom[9],rom[8]} = 32'b00000000000000000000000000010011;
        {rom[15],rom[14],rom[13],rom[12]} = 32'b00000000010100101000001100110011;
        {rom[19],rom[18],rom[17],rom[16]} = 32'b00000000000000000000000000010011;
        {rom[23],rom[22],rom[21],rom[20]} = 32'b00000000000000000000000000010011;
        {rom[27],rom[26],rom[25],rom[24]} = 32'b01000000011000000000001110110011;
        {rom[31],rom[30],rom[29],rom[28]} = 32'b00000000011000101111111000110011;
        {rom[35],rom[34],rom[33],rom[32]} = 32'b00000000001000000000111000010011;
        {rom[39],rom[38],rom[37],rom[36]} = 32'b00000000000000000000000000010011;
        {rom[43],rom[42],rom[41],rom[40]} = 32'b00000000000000000000000000010011;
        {rom[47],rom[46],rom[45],rom[44]} = 32'b00000001110000110001001100110011;
        {rom[51],rom[50],rom[49],rom[48]} = 32'b00000000000000000000000000010011;
        {rom[55],rom[54],rom[53],rom[52]} = 32'b00000000000000000000000000010011;
        {rom[59],rom[58],rom[57],rom[56]} = 32'b00000000011000111110001110110011;
        {rom[63],rom[62],rom[61],rom[60]} = 32'b00000000000000000000000000010011;
        {rom[67],rom[66],rom[65],rom[64]} = 32'b00000000000000000000000000010011;
        {rom[71],rom[70],rom[69],rom[68]} = 32'b01110011001000111111111010010011;
        {rom[75],rom[74],rom[73],rom[72]} = 32'b00000000000000000000000000010011;
        {rom[79],rom[78],rom[77],rom[76]} = 32'b00000000000000000000000000010011;
        {rom[83],rom[82],rom[81],rom[80]} = 32'b00000000010111101101111010010011;
        {rom[87],rom[86],rom[85],rom[84]} = 32'b00000000000000000000000000010011;
        {rom[91],rom[90],rom[89],rom[88]} = 32'b00000000000000000000000000010011;
        {rom[95],rom[94],rom[93],rom[92]} = 32'b00000001110000111101001110110011;
        {rom[99],rom[98],rom[97],rom[96]} = 32'b00000000000000000000000000010011;
        {rom[103],rom[102],rom[101],rom[100]} = 32'b00000000000000000000000000010011;
        {rom[107],rom[106],rom[105],rom[104]} = 32'b00000001000000111001001110010011;
        {rom[111],rom[110],rom[109],rom[108]} = 32'b00000000000000000000000000010011;
        {rom[115],rom[114],rom[113],rom[112]} = 32'b00000000000000000000000000010011;
        {rom[119],rom[118],rom[117],rom[116]} = 32'b01000001110000111101001110110011;
        {rom[123],rom[122],rom[121],rom[120]} = 32'b00000000011000101001100001100011;////////////
        {rom[127],rom[126],rom[125],rom[124]} = 32'b00000000000000000000000000010011;
        {rom[131],rom[130],rom[129],rom[128]} = 32'b00000000000000000000000000010011;
        {rom[135],rom[134],rom[133],rom[132]} = 32'b00000000000000000000001110110011;
        {rom[139],rom[138],rom[137],rom[136]} = 32'b00000010000000111000100001100011;
        {rom[143],rom[142],rom[141],rom[140]} = 32'b00000000000000000000000000010011;
        {rom[147],rom[146],rom[145],rom[144]} = 32'b00000000000000000000000000010011;
        {rom[151],rom[150],rom[149],rom[148]} = 32'b00000011110100111101001001100011;
        {rom[155],rom[154],rom[153],rom[152]} = 32'b00000000000000000000000000010011;
        {rom[159],rom[158],rom[157],rom[156]} = 32'b00000000000000000000000000010011;
        {rom[163],rom[162],rom[161],rom[160]} = 32'b00000000000000111000001010110011;
        {rom[167],rom[166],rom[165],rom[164]} = 32'b00000000000000000000000000010011;
        {rom[171],rom[170],rom[169],rom[168]} = 32'b00000000000000000000000000010011;
        {rom[175],rom[174],rom[173],rom[172]} = 32'b00000001110100111100100001100011;
        {rom[179],rom[178],rom[177],rom[176]} = 32'b00000000000000000000000000010011;
        {rom[183],rom[182],rom[181],rom[180]} = 32'b00000000000000000000000000010011;
        {rom[187],rom[186],rom[185],rom[184]} = 32'b00000000000000000000001010110011;
        {rom[191],rom[190],rom[189],rom[188]} = 32'b00000000010100111001110001100011;
        {rom[195],rom[194],rom[193],rom[192]} = 32'b00000000000000000000000000010011;
        {rom[199],rom[198],rom[197],rom[196]} = 32'b00000000000000000000000000010011;
        {rom[203],rom[202],rom[201],rom[200]} = 32'b00000000010100111000100001100011;
        {rom[207],rom[206],rom[205],rom[204]} = 32'b00000000000000000000000000010011;
        {rom[211],rom[210],rom[209],rom[208]} = 32'b00000000000000000000000000010011;
        {rom[215],rom[214],rom[213],rom[212]} = 32'b00000000000000000000001100110011;
        {rom[219],rom[218],rom[217],rom[216]} = 32'b00000001110100110100110001100011;
        {rom[223],rom[222],rom[221],rom[220]} = 32'b00000000000000000000000000010011;
        {rom[227],rom[226],rom[225],rom[224]} = 32'b00000000000000000000000000010011;
        {rom[231],rom[230],rom[229],rom[228]} = 32'b00000001110000110101100001100011;
        {rom[235],rom[234],rom[233],rom[232]} = 32'b00000000000000000000000000010011;
        {rom[239],rom[238],rom[237],rom[236]} = 32'b00000000000000000000000000010011;
        {rom[243],rom[242],rom[241],rom[240]} = 32'b00000000000000000000111000110011;
        {rom[247],rom[246],rom[245],rom[244]} = 32'b00000000000000000000111010110011;
        {rom[251],rom[250],rom[249],rom[248]} = 32'b00000001100000000000000011101111;
        {rom[255],rom[254],rom[253],rom[252]} = 32'b00000000000000000000000000010011;
        {rom[259],rom[258],rom[257],rom[256]} = 32'b00000000000000000000000000010011;
        {rom[263],rom[262],rom[261],rom[260]} = 32'b00000010011100101000100001100011;
        {rom[267],rom[266],rom[265],rom[264]} = 32'b00000000000000000000000000010011;
        {rom[271],rom[270],rom[269],rom[268]} = 32'b00000000000000000000000000010011;
        {rom[275],rom[274],rom[273],rom[272]} = 32'b00000000010100010010000000100011;
        {rom[279],rom[278],rom[277],rom[276]} = 32'b00000000011000010000001000100011;
        {rom[283],rom[282],rom[281],rom[280]} = 32'b00000000000000010010111010000011;
        {rom[287],rom[286],rom[285],rom[284]} = 32'b00000000010000010000111010000011;
        {rom[291],rom[290],rom[289],rom[288]} = 32'b00000000010000010100111010000011;
        {rom[295],rom[294],rom[293],rom[292]} = 32'b00000000000000001000000001100111;
        {rom[299],rom[298],rom[297],rom[296]} = 32'b00000000000000000000000000010011;
        {rom[303],rom[302],rom[301],rom[300]} = 32'b00000000000000000000000000010011;
        {rom[307],rom[306],rom[305],rom[304]} = 32'b00000000000000000000000010110011;
        {rom[311],rom[310],rom[309],rom[308]} = 32'b00000000000000000000001110110011;
    end
    
    always@(*)
        instruction = {rom[cur_pc + 3], rom[cur_pc + 2], rom[cur_pc + 1], rom[cur_pc]};
            
endmodule

